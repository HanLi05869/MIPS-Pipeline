`timescale 1ns / 1ps

module IM(
		input[11:2] addr,
		output reg[31:0] IS
	);
	reg[31:0] im[1023:0];
	integer i;
	always @addr
	begin
		IS = im[addr];
	end

    /*
    initial begin
        $readmemh("TESTCODE.txt", im, 0, 1023);
    end
    */
	//test
	initial
	begin
		for(i = 0; i < 1024; i += 1) 
			im[i] = 0;

		/*im[0] = 32'b10001100000000010000000000000100;
		im[1] = 32'b10001100000000100000000000001000;
		im[2] = 32'b00000000001000100001100000100001;
		im[3] = 32'b00000000010000110010000000100001;
		im[4] = 32'b00000000011001000010100000100001;
		im[5] = 32'b00000000100001010011000000100001;
		*/
		/*im[0] = 32'b00100000101001010000000000000001;//addi
		im[1] = 32'b10101100000001010000000000000100;//sw
		im[2] = 32'b10101100000001010000000000001000;//sw
		im[3] = 32'b00000000101001010011000000100001;//addu
		im[4] = 32'b10101100000001100000000000001100;//sw
		im[5] = 32'b10101100000001100000000000010000;//sw
		im[6] = 32'b00110100111001110000000000000100;//ori
		im[7] = 32'b10001100111010000000000000000100;//lw
		im[8] = 32'b00000000111001100100100000100011;//subu
		im[9] = 32'b00010001001001100000000000000001;//beq
		im[10] = 32'b00000001001010010100100000100001;//addu
		im[11] = 32'b00000000111010010101000000101010;//slt
		im[12] = 32'b00010001010000000000000000000001;//beq
		im[13] = 32'b00000001001010010100100000100001;//addu
		im[14] = 32'b00001000000000000000110000010001;//j
		im[15] = 32'b00000001001010010110000000100001;//addu
		im[16] = 32'b00000011111000000000000000001000;//jr
		im[17] = 32'b00111100000010110000000000000001;//lui
		im[18] = 32'b00001100000000000000110000001111;//jal
		im[19] = 32'b00000001100010000110100000100011;//subu*/

	
		
		im[0] = 32'b00110100101001010000000000000001;
        im[1] = 32'b00000000101001010110100000100001;
        im[2] = 32'b00100000110001100000000000000100;
        im[3] = 32'b10101100110001100000000000000000;
        im[4] = 32'b10001100000001110000000000000100;
        im[5] = 32'b00000000101001110100000000101010;
        im[6] = 32'b00010001000001010000000000000001;
        im[7] = 32'b00000001000010000100000000100011;
        im[8] = 32'b00000000111001010100100000100011;
        im[9] = 32'b00001000000000000000110000001100;
        im[10] = 32'b00000000110010100101100000100011;
        im[11] = 32'b00000011111000000000000000001000;
        im[12] = 32'b00111100000010100000000000000001;
        im[13] = 32'b00001100000000000000110000001010;
        im[14] = 32'b00110101100011000000000000001100;

/**/
	end
    
endmodule